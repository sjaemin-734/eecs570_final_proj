SET_CLAUSE_DATABASE(0, 55'b0000000000000000000000000000000000000000000000000000000);
SET_CLAUSE_DATABASE(1, 55'b1110000011000000001000000010000000011000000000000000000);
SET_CLAUSE_DATABASE(2, 55'b1110000111000000001000000010000000011000000000000000000);
SET_CLAUSE_DATABASE(3, 55'b1110001011000000001000000010000000011000000000000000000);
SET_CLAUSE_DATABASE(4, 55'b1110001111000000001000000010000000011000000000000000000);
SET_CLAUSE_DATABASE(5, 55'b1110010011000000001000000010000000011000000000000000000);
SET_CLAUSE_DATABASE(6, 55'b1110010111000000001000000010000000011000000000000000000);
SET_CLAUSE_DATABASE(7, 55'b1110011011000000001000000010000000011000000000000000000);
SET_CLAUSE_DATABASE(8, 55'b1110011111000000001000000010000000011000000000000000000);