`ifndef __SYS_DEFS_SVH__
`define __SYS_DEFS_SVH__

`define MAX_VARS 512
`define MAX_CLAUSES 1024


`endif // __SYS_DEFS_SVH__