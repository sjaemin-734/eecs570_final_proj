`ifndef __SYS_DEFS_SVH__
`define __SYS_DEFS_SVH__

`define MAX_VARS 512
`define MAX_VARS_BITS $clog2(MAX_VARS)
`define MAX_CLAUSES 1024
`define MAX_CLAUSES_BITS $clog2(MAX_CLAUSES)
`define VAR_PER_CLAUSE 5


`endif // __SYS_DEFS_SVH__